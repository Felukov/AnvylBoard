library IEEE;
library UNISIM;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use UNISIM.VComponents.all;
use ieee.math_real.all;

entity vid_mem_ctrl is
    port (
        clk   : in std_logic;
        reset : in std_logic

    );
end entity vid_mem_ctrl;

architecture rtl of vid_mem_ctrl is

begin



end architecture;