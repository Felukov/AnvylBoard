library ieee;
library unisim;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use unisim.vcomponents.all;

entity vid_mem_glyph is
    port (
        clk         : in std_logic;
        glyph_addr  : in std_logic_vector(10 downto 0);
        glyph_line  : out std_logic_vector(39 downto 0)
    );
end entity vid_mem_glyph;

architecture rtl of vid_mem_glyph is

    --12x8 matrix
	type rom_type is array (0 to 34*31-1) of std_logic_vector(39 downto 0);

    signal rom : rom_type := (
        --0
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000011111111111111111111111100000000",
        "0000000111111111111111111111111110000000",
        "0000001111111111111111111111111111000000",
        "0000001110000000000000000000111111000000",
        "0000001110000000000000000001110111000000",
        "0000001110000000000000000011100111000000",
        "0000001110000000000000000111000111000000",
        "0000001110000000000000001110000111000000",
        "0000001110000000000000011100000111000000",
        "0000001110000000000000111000000111000000",
        "0000001110000000000001110000000111000000",
        "0000001110000000000011100000000111000000",
        "0000001110000000000111000000000111000000",
        "0000001110000000001110000000000111000000",
        "0000001110000000011100000000000111000000",
        "0000001110000000111000000000000111000000",
        "0000001110000001110000000000000111000000",
        "0000001110000011100000000000000111000000",
        "0000001110000111000000000000000111000000",
        "0000001110001110000000000000000111000000",
        "0000001110011100000000000000000111000000",
        "0000001110111000000000000000000111000000",
        "0000001111110000000000000000000111000000",
        "0000001111111111111111111111111111000000",
        "0000000111111111111111111111111110000000",
        "0000000011111111111111111111111100000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        --1
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000011110000000000000000000",
        "0000000000000000111110000000000000000000",
        "0000000000000001111110000000000000000000",
        "0000000000000011101110000000000000000000",
        "0000000000000111001110000000000000000000",
        "0000000000001110001110000000000000000000",
        "0000000000011100001110000000000000000000",
        "0000000000111000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        --2
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000111111111111111111110000000000",
        "0000000011111111111111111111111100000000",
        "0000001111111111111111111111111110000000",
        "0000001111100000000000000000011111000000",
        "0000001111000000000000000000001111000000",
        "0000001110000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000001111000000",
        "0000000000000000000000000001111110000000",
        "0000000000000000000000000111111000000000",
        "0000000000000000000001111111100000000000",
        "0000000000000000011111111100000000000000",
        "0000000000000111111111000000000000000000",
        "0000000000111111110000000000000000000000",
        "0000000011111110000000000000000000000000",
        "0000001111110000000000000000000000000000",
        "0000001111000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000001111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        --3
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000011111111111111111111111100000000",
        "0000000111111111111111111111111110000000",
        "0000001111111111111111111111111111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000001111000000",
        "0000000000000000000000000000111111000000",
        "0000000000000000111111111111111110000000",
        "0000000000000011111111111111111000000000",
        "0000000000000001111111111111111110000000",
        "0000000000000000000000000000001111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001111000000000000000000001111000000",
        "0000001111110000000000000000111111000000",
        "0000000111111111111111111111111110000000",
        "0000000011111111111111111111111000000000",
        "0000000000111111111111111111100000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        --3
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000111000000000111000000",
        "0000000000000000001110000000000111000000",
        "0000000000000000011100000000000111000000",
        "0000000000000000111000000000000111000000",
        "0000000000000001110000000000000111000000",
        "0000000000000011100000000000000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000001110000000000000000111000000",
        "0000000000011100000000000000000111000000",
        "0000000000111000000000000000000111000000",
        "0000000001110000000000000000000111000000",
        "0000000011100000000000000000000111000000",
        "0000000111000000000000000000000111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        --5
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110111111111111111111110000000000",
        "0000001111111111111111111111111000000000",
        "0000001111111111111111111111111110000000",
        "0000001111000000000000000000111111000000",
        "0000001110000000000000000000001111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000001110000000000000000000001111000000",
        "0000001111000000000000000000111111000000",
        "0000001111111111111111111111111111000000",
        "0000000111111111111111111111111110000000",
        "0000000001111111111111111111110000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --6
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000011111111111111111111111110000000",
        "0000000111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001111000000000000000000000111000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110011111111111111111110000000000",
        "0000001111111111111111111111111000000000",
        "0000001111111111111111111111111110000000",
        "0000001111100000000000000000011111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001111100000000000000000011111000000",
        "0000001111111111111111111111111111000000",
        "0000000111111111111111111111111110000000",
        "0000000011111111111111111111111100000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --7
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000111111111111111111111111110000000",
        "0000000111111111111111111111111110000000",
        "0000000111111111111111111111111110000000",
        "0000000111000000000000000000011100000000",
        "0000000000000000000000000000111000000000",
        "0000000000000000000000000000111000000000",
        "0000000000000000000000000001110000000000",
        "0000000000000000000000000001110000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000111000000000000",
        "0000000000000000000000000111000000000000",
        "0000000000000000000000001110000000000000",
        "0000000000000000000000001110000000000000",
        "0000000000000000000000011100000000000000",
        "0000000000000000000000011100000000000000",
        "0000000000000000000000111000000000000000",
        "0000000000000000000000111000000000000000",
        "0000000000000000000001110000000000000000",
        "0000000000000000000001110000000000000000",
        "0000000000000000000011100000000000000000",
        "0000000000000000000011100000000000000000",
        "0000000000000000000111000000000000000000",
        "0000000000000000000111000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --8
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000111111111111111111110000000000",
        "0000000111111111111111111111111110000000",
        "0000001111111111111111111111111111000000",
        "0000001111100000000000000000011111000000",
        "0000001111000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001111000000000000000000001111000000",
        "0000000111110000000000000000111110000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000111111111111111111111111110000000",
        "0000001111000000000000000000001111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001111000000000000000000001111000000",
        "0000001111111111111111111111111111000000",
        "0000000111111111111111111111111110000000",
        "0000000011111111111111111111111100000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --9
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000111111111111111111110000000000",
        "0000000111111111111111111111111110000000",
        "0000001111111111111111111111111111000000",
        "0000001111100000000000000000011111000000",
        "0000001111000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001111000000000000000000000111000000",
        "0000000111110000000000000000000111000000",
        "0000000011111111111111111111111111000000",
        "0000000000111111111111111111111111000000",
        "0000000000011111111111111111111111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000000000000000000000000000000111000000",
        "0000001111000000000000000000001111000000",
        "0000001111111111111111111111111111000000",
        "0000000111111111111111111111111110000000",
        "0000000011111111111111111111111100000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --A
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000001110000000000000000000",
        "0000000000000000011111000000000000000000",
        "0000000000000000111111100000000000000000",
        "0000000000000000111111100000000000000000",
        "0000000000000001110001110000000000000000",
        "0000000000000001110001110000000000000000",
        "0000000000000011100000111000000000000000",
        "0000000000000011100000111000000000000000",
        "0000000000000111000000011100000000000000",
        "0000000000000111000000011100000000000000",
        "0000000000001110000000001110000000000000",
        "0000000000001110000000001110000000000000",
        "0000000000011100000000000111000000000000",
        "0000000000011111111111111111000000000000",
        "0000000000111111111111111111100000000000",
        "0000000000111000000000000011100000000000",
        "0000000001110000000000000001110000000000",
        "0000000001110000000000000001110000000000",
        "0000000011100000000000000000111000000000",
        "0000000011100000000000000000111000000000",
        "0000000111000000000000000000011100000000",
        "0000000111000000000000000000011100000000",
        "0000001110000000000000000000001110000000",
        "0000001110000000000000000000001110000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --B
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000001111111111111111111111110000000000",
        "0000001111111111111111111111111110000000",
        "0000001111111111111111111111111111000000",
        "0000001110000000000000000000011111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000001111000000",
        "0000001110000000000000000000111110000000",
        "0000001111111111111111111111111000000000",
        "0000001111111111111111111111111000000000",
        "0000001111111111111111111111111110000000",
        "0000001110000000000000000000001111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000001111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111110000000",
        "0000001111111111111111111111111100000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --C
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000111111111111111111110000000000",
        "0000000111111111111111111111111110000000",
        "0000001111111111111111111111111111000000",
        "0000001111100000000000000000011111000000",
        "0000001111000000000000000000000111000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000111000000",
        "0000001111000000000000000000001111000000",
        "0000001111111111111111111111111111000000",
        "0000000111111111111111111111111110000000",
        "0000000011111111111111111111111100000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --D
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000001111111111111111111111110000000000",
        "0000001111111111111111111111111110000000",
        "0000001111111111111111111111111111000000",
        "0000001110000000000000000000011111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000000111000000",
        "0000001110000000000000000000001111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111110000000",
        "0000001111111111111111111111111100000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --E
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001110000000000000000000011111000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001111111111111111111111111000000000",
        "0000001111111111111111111111111000000000",
        "0000001111111111111111111111111000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000001111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --F
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001111111111111111111111111111000000",
        "0000001110000000000000000000011111000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001111111111111111111111111000000000",
        "0000001111111111111111111111111000000000",
        "0000001111111111111111111111111000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000001110000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --+
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        -- -
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --*
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000001110000001111000000111000000000",
        "0000000001110000001111000000111000000000",
        "0000000001110000001111000000111000000000",
        "0000000000001110001111000111000000000000",
        "0000000000001110001111000111000000000000",
        "0000000000001110001111000111000000000000",
        "0000000000000001111111111000000000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000000000001111111111000000000000000",
        "0000000000001110001111000111000000000000",
        "0000000000001110001111000111000000000000",
        "0000000000001110001111000111000000000000",
        "0000000001110000001111000000111000000000",
        "0000000001110000001111000000111000000000",
        "0000000001110000001111000000111000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --/
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --AND
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011100000000000000111000000000000000",
        "0000011100000000000000111000000000000000",
        "0000011100000111111111111111111111000000",
        "0000011100000111111111111111111111000000",
        "0000011100000111111111111111111111000000",
        "0000011100000111111111111100000111000000",
        "0000011100000111111111111100000111000000",
        "0000011100000111111111111100000111000000",
        "0000011111111111111111111100000111000000",
        "0000011111111111111111111100000111000000",
        "0000011111111111111111111100000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --OR
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111111111111000000",
        "0000011111111111111111111111111111000000",
        "0000011111111111111111111111111111000000",
        "0000011111111111111111111111111111000000",
        "0000011111111111111111111111111111000000",
        "0000011111111111111111111111111111000000",
        "0000011111111111111111111111111111000000",
        "0000011111111111111111111111111111000000",
        "0000011111111111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --AND
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011111111111111111111000000000000000",
        "0000011100000000000000111000000000000000",
        "0000011100000000000000111000000000000000",
        "0000011100000111111111111111111111000000",
        "0000011100000111111111111111111111000000",
        "0000011100000111111111111111111111000000",
        "0000011100000111000000111100000111000000",
        "0000011100000111000000111100000111000000",
        "0000011100000111000000111100000111000000",
        "0000011111111111111111111100000111000000",
        "0000011111111111111111111100000111000000",
        "0000011111111111111111111100000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000000111000000000000000111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000111111111111111111111000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --/
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",


        --1
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000111100000000000",
        "0000000000000000000000001111100000000000",
        "0000000000000000000000011111100000000000",
        "0000000000000000000000111011100000000000",
        "0000000000000000000001110011100000000000",
        "0000000000000000000011100011100000000000",
        "0000000000000000000111000011100000000000",
        "0000000000000000001110000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000001111111111111100000011100000000000",
        "0000001111111111111100000011100000000000",
        "0000001111111111111100000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000000000011100000000000",
        "0000000000000000000001111111111111000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --shl
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000001000000000000010000000",
        "0000000000000000011000000000000110000000",
        "0000000000000000111000000000001110000000",
        "0000000000000001111000000000011110000000",
        "0000000000000011111000000000111110000000",
        "0000000000000111111000000001111110000000",
        "0000000000001111111000000011111110000000",
        "0000000000011111111000000111111110000000",
        "0000000000111111111000001111111110000000",
        "0000000001111111111000011111111110000000",
        "0000000011111111111000111111111110000000",
        "0000000111111111111001111111111110000000",
        "0000001111111111111011111111111110000000",
        "0000000111111111111001111111111110000000",
        "0000000011111111111000111111111110000000",
        "0000000001111111111000011111111110000000",
        "0000000000111111111000001111111110000000",
        "0000000000011111111000000111111110000000",
        "0000000000001111111000000011111110000000",
        "0000000000000111111000000001111110000000",
        "0000000000000011111000000000111110000000",
        "0000000000000001111000000000011110000000",
        "0000000000000000111000000000001110000000",
        "0000000000000000011000000000000110000000",
        "0000000000000000001000000000000010000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --shl
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000010000000000001000000000000000000",
        "0000000011000000000001100000000000000000",
        "0000000011100000000001110000000000000000",
        "0000000011110000000001111000000000000000",
        "0000000011111000000001111100000000000000",
        "0000000011111100000001111110000000000000",
        "0000000011111110000001111111000000000000",
        "0000000011111111000001111111100000000000",
        "0000000011111111100001111111110000000000",
        "0000000011111111110001111111111000000000",
        "0000000011111111111001111111111100000000",
        "0000000011111111111101111111111110000000",
        "0000000011111111111111111111111111000000",
        "0000000011111111111101111111111110000000",
        "0000000011111111111001111111111100000000",
        "0000000011111111110001111111111000000000",
        "0000000011111111100001111111110000000000",
        "0000000011111111000001111111100000000000",
        "0000000011111110000001111111000000000000",
        "0000000011111100000001111110000000000000",
        "0000000011111000000001111100000000000000",
        "0000000011110000000001111000000000000000",
        "0000000011100000000001110000000000000000",
        "0000000011000000000001100000000000000000",
        "0000000010000000000001000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --/
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000001111111111111111111111000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --back
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000100000000000000000000",
        "0000000000000000001100000000000000000000",
        "0000000000000000011100000000000000000000",
        "0000000000000000111100000000000000000000",
        "0000000000000001111100000000000000000000",
        "0000000000000011111100000000000000000000",
        "0000000000000111111100000000000000000000",
        "0000000000001111111100000000000000000000",
        "0000000000011111111100000000000000000000",
        "0000000000111111111100000000000000000000",
        "0000000001111111111111111111111111000000",
        "0000000011111111111111111111111111000000",
        "0000000111111111111111111111111111000000",
        "0000000011111111111111111111111111000000",
        "0000000001111111111111111111111111000000",
        "0000000000111111111100000000000000000000",
        "0000000000011111111100000000000000000000",
        "0000000000001111111100000000000000000000",
        "0000000000000111111100000000000000000000",
        "0000000000000011111100000000000000000000",
        "0000000000000001111100000000000000000000",
        "0000000000000000111100000000000000000000",
        "0000000000000000011100000000000000000000",
        "0000000000000000001100000000000000000000",
        "0000000000000000000100000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --null
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",

        --/
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000001111000000000000000000000000000",
        "0000000001111000000000000011110000000000",
        "0000000001111000000000000011110000000000",
        "0000000000000000000000000111110000000000",
        "0000000000000000000000111110000000000000",
        "0000000000000000000000111100000000000000",
        "0000000000000000000001111100000000000000",
        "0000000000000000001111100000000000000000",
        "0000000000000000001111000000000000000000",
        "0000000000000000011111000000000000000000",
        "0000000000000011111000000000000000000000",
        "0000000000000011110000000000000000000000",
        "0000000000000111110000000000000000000000",
        "0000000000111110000000000000000000000000",
        "0000000000111100000000000001111000000000",
        "0000000000111100000000000001111000000000",
        "0000000000000000000000000001111000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000"
    );


begin

	fetch_line_process: process (clk) begin
		if rising_edge(clk) then
			-- Read from Rom
			glyph_line <= rom(to_integer(unsigned(glyph_addr)));
		end if;
	end process;

end architecture;