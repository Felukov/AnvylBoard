library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

entity cpu_ctrl is

    port (
        cpu_clk         : in std_logic
    );

end cpu_ctrl;

architecture Behavioral of cpu_ctrl is


begin

end Behavioral;
