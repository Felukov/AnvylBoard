library ieee;
library unisim;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use unisim.vcomponents.all;

entity oled_char_lib is
    port (
        clk   : in std_logic;
        addra : in std_logic_vector(10 downto 0); --first 8 bits is the ascii value of the character the last 3 bits are the parts of the char
        douta : out std_logic_vector(7 downto 0) --data byte out

    );
end entity oled_char_lib;

architecture rtl of oled_char_lib is
    type rom_type_t is array (0 to 1023) of std_logic_vector(7 downto 0);
    signal rom : rom_type_t := (
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01011111",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000011",
        "00000000",
        "00000011",
        "00000000",
        "00000000",
        "00000000",
        "01100100",
        "00111100",
        "00100110",
        "01100100",
        "00111100",
        "00100110",
        "00100100",
        "00000000",
        "00100110",
        "01001001",
        "01001001",
        "01111111",
        "01001001",
        "01001001",
        "00110010",
        "00000000",
        "01000010",
        "00100101",
        "00010010",
        "00001000",
        "00100100",
        "01010010",
        "00100001",
        "00000000",
        "00100000",
        "01010000",
        "01001110",
        "01010101",
        "00100010",
        "01011000",
        "00101000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000011",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00011100",
        "00100010",
        "01000001",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000001",
        "00100010",
        "00011100",
        "00000000",
        "00000000",
        "00000000",
        "00010101",
        "00010101",
        "00001110",
        "00001110",
        "00010101",
        "00010101",
        "00000000",
        "00000000",
        "00001000",
        "00001000",
        "00111110",
        "00001000",
        "00001000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01010000",
        "00110000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00001000",
        "00001000",
        "00001000",
        "00001000",
        "00001000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000000",
        "00100000",
        "00010000",
        "00001000",
        "00000100",
        "00000010",
        "00000001",
        "00000000",
        "00000000",
        "00111110",
        "01000001",
        "01000001",
        "01000001",
        "00111110",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000001",
        "01111111",
        "01000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000010",
        "01100001",
        "01010001",
        "01001001",
        "01101110",
        "00000000",
        "00000000",
        "00000000",
        "00100010",
        "01000001",
        "01001001",
        "01001001",
        "00110110",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00010100",
        "00010010",
        "01111111",
        "00010000",
        "00000000",
        "00000000",
        "00000000",
        "00100111",
        "01001001",
        "01001001",
        "01001001",
        "01110001",
        "00000000",
        "00000000",
        "00000000",
        "00111100",
        "01001010",
        "01001001",
        "01001000",
        "01110000",
        "00000000",
        "00000000",
        "00000000",
        "01000011",
        "00100001",
        "00010001",
        "00001101",
        "00000011",
        "00000000",
        "00000000",
        "00000000",
        "00110110",
        "01001001",
        "01001001",
        "01001001",
        "00110110",
        "00000000",
        "00000000",
        "00000000",
        "00000110",
        "00001001",
        "01001001",
        "00101001",
        "00011110",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00010010",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01010010",
        "00110000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00001000",
        "00010100",
        "00010100",
        "00100010",
        "00000000",
        "00000000",
        "00000000",
        "00010100",
        "00010100",
        "00010100",
        "00010100",
        "00010100",
        "00010100",
        "00000000",
        "00000000",
        "00000000",
        "00100010",
        "00010100",
        "00010100",
        "00001000",
        "00000000",
        "00000000",
        "00000000",
        "00000010",
        "00000001",
        "01011001",
        "00000101",
        "00000010",
        "00000000",
        "00000000",
        "00111110",
        "01000001",
        "01011101",
        "01010101",
        "01001101",
        "01010001",
        "00101110",
        "00000000",
        "01000000",
        "01111100",
        "01001010",
        "00001001",
        "01001010",
        "01111100",
        "01000000",
        "00000000",
        "01000001",
        "01111111",
        "01001001",
        "01001001",
        "01001001",
        "01001001",
        "00110110",
        "00000000",
        "00011100",
        "00100010",
        "01000001",
        "01000001",
        "01000001",
        "01000001",
        "00100010",
        "00000000",
        "01000001",
        "01111111",
        "01000001",
        "01000001",
        "01000001",
        "00100010",
        "00011100",
        "00000000",
        "01000001",
        "01111111",
        "01001001",
        "01001001",
        "01011101",
        "01000001",
        "01100011",
        "00000000",
        "01000001",
        "01111111",
        "01001001",
        "00001001",
        "00011101",
        "00000001",
        "00000011",
        "00000000",
        "00011100",
        "00100010",
        "01000001",
        "01001001",
        "01001001",
        "00111010",
        "00001000",
        "00000000",
        "01000001",
        "01111111",
        "00001000",
        "00001000",
        "00001000",
        "01111111",
        "01000001",
        "00000000",
        "00000000",
        "01000001",
        "01000001",
        "01111111",
        "01000001",
        "01000001",
        "00000000",
        "00000000",
        "00110000",
        "01000000",
        "01000001",
        "01000001",
        "00111111",
        "00000001",
        "00000001",
        "00000000",
        "01000001",
        "01111111",
        "00001000",
        "00001100",
        "00010010",
        "01100001",
        "01000001",
        "00000000",
        "01000001",
        "01111111",
        "01000001",
        "01000000",
        "01000000",
        "01000000",
        "01100000",
        "00000000",
        "01000001",
        "01111111",
        "01000010",
        "00001100",
        "01000010",
        "01111111",
        "01000001",
        "00000000",
        "01000001",
        "01111111",
        "01000010",
        "00001100",
        "00010001",
        "01111111",
        "00000001",
        "00000000",
        "00011100",
        "00100010",
        "01000001",
        "01000001",
        "01000001",
        "00100010",
        "00011100",
        "00000000",
        "01000001",
        "01111111",
        "01001001",
        "00001001",
        "00001001",
        "00001001",
        "00000110",
        "00000000",
        "00001100",
        "00010010",
        "00100001",
        "00100001",
        "01100001",
        "01010010",
        "01001100",
        "00000000",
        "01000001",
        "01111111",
        "00001001",
        "00001001",
        "00011001",
        "01101001",
        "01000110",
        "00000000",
        "01100110",
        "01001001",
        "01001001",
        "01001001",
        "01001001",
        "01001001",
        "00110011",
        "00000000",
        "00000011",
        "00000001",
        "01000001",
        "01111111",
        "01000001",
        "00000001",
        "00000011",
        "00000000",
        "00000001",
        "00111111",
        "01000001",
        "01000000",
        "01000001",
        "00111111",
        "00000001",
        "00000000",
        "00000001",
        "00001111",
        "00110001",
        "01000000",
        "00110001",
        "00001111",
        "00000001",
        "00000000",
        "00000001",
        "00011111",
        "01100001",
        "00010100",
        "01100001",
        "00011111",
        "00000001",
        "00000000",
        "01000001",
        "01000001",
        "00110110",
        "00001000",
        "00110110",
        "01000001",
        "01000001",
        "00000000",
        "00000001",
        "00000011",
        "01000100",
        "01111000",
        "01000100",
        "00000011",
        "00000001",
        "00000000",
        "01000011",
        "01100001",
        "01010001",
        "01001001",
        "01000101",
        "01000011",
        "01100001",
        "00000000",
        "00000000",
        "00000000",
        "01111111",
        "01000001",
        "01000001",
        "00000000",
        "00000000",
        "00000000",
        "00000001",
        "00000010",
        "00000100",
        "00001000",
        "00010000",
        "00100000",
        "01000000",
        "00000000",
        "00000000",
        "00000000",
        "01000001",
        "01000001",
        "01111111",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000100",
        "00000010",
        "00000001",
        "00000001",
        "00000010",
        "00000100",
        "00000000",
        "00000000",
        "01000000",
        "01000000",
        "01000000",
        "01000000",
        "01000000",
        "01000000",
        "00000000",
        "00000000",
        "00000001",
        "00000010",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00110100",
        "01001010",
        "01001010",
        "01001010",
        "00111100",
        "01000000",
        "00000000",
        "00000000",
        "01000001",
        "00111111",
        "01001000",
        "01001000",
        "01001000",
        "00110000",
        "00000000",
        "00000000",
        "00111100",
        "01000010",
        "01000010",
        "01000010",
        "00100100",
        "00000000",
        "00000000",
        "00000000",
        "00110000",
        "01001000",
        "01001000",
        "01001001",
        "00111111",
        "01000000",
        "00000000",
        "00000000",
        "00111100",
        "01001010",
        "01001010",
        "01001010",
        "00101100",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01001000",
        "01111110",
        "01001001",
        "00001001",
        "00000000",
        "00000000",
        "00000000",
        "00100110",
        "01001001",
        "01001001",
        "01001001",
        "00111111",
        "00000001",
        "00000000",
        "01000001",
        "01111111",
        "01001000",
        "00000100",
        "01000100",
        "01111000",
        "01000000",
        "00000000",
        "00000000",
        "00000000",
        "01000100",
        "01111101",
        "01000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000000",
        "01000100",
        "00111101",
        "00000000",
        "00000000",
        "00000000",
        "01000001",
        "01111111",
        "00010000",
        "00011000",
        "00100100",
        "01000010",
        "01000010",
        "00000000",
        "00000000",
        "01000000",
        "01000001",
        "01111111",
        "01000000",
        "01000000",
        "00000000",
        "00000000",
        "01000010",
        "01111110",
        "00000010",
        "01111100",
        "00000010",
        "01111110",
        "01000000",
        "00000000",
        "01000010",
        "01111110",
        "01000100",
        "00000010",
        "01000010",
        "01111100",
        "01000000",
        "00000000",
        "00000000",
        "00111100",
        "01000010",
        "01000010",
        "01000010",
        "00111100",
        "00000000",
        "00000000",
        "00000000",
        "01000001",
        "01111111",
        "01001001",
        "00001001",
        "00001001",
        "00000110",
        "00000000",
        "00000000",
        "00000110",
        "00001001",
        "00001001",
        "01001001",
        "01111111",
        "01000001",
        "00000000",
        "00000000",
        "01000010",
        "01111110",
        "01000100",
        "00000010",
        "00000010",
        "00000100",
        "00000000",
        "00000000",
        "01100100",
        "01001010",
        "01001010",
        "01001010",
        "00110110",
        "00000000",
        "00000000",
        "00000000",
        "00000100",
        "00111111",
        "01000100",
        "01000100",
        "00100000",
        "00000000",
        "00000000",
        "00000000",
        "00000010",
        "00111110",
        "01000000",
        "01000000",
        "00100010",
        "01111110",
        "01000000",
        "00000010",
        "00001110",
        "00110010",
        "01000000",
        "00110010",
        "00001110",
        "00000010",
        "00000000",
        "00000010",
        "00011110",
        "01100010",
        "00011000",
        "01100010",
        "00011110",
        "00000010",
        "00000000",
        "01000010",
        "01100010",
        "00010100",
        "00001000",
        "00010100",
        "01100010",
        "01000010",
        "00000000",
        "00000001",
        "01000011",
        "01000101",
        "00111000",
        "00000101",
        "00000011",
        "00000001",
        "00000000",
        "00000000",
        "01000110",
        "01100010",
        "01010010",
        "01001010",
        "01000110",
        "01100010",
        "00000000",
        "00000000",
        "00000000",
        "00001000",
        "00110110",
        "01000001",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01111111",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "00000000",
        "01000001",
        "00110110",
        "00001000",
        "00000000",
        "00000000",
        "00000000",
        "00011000",
        "00001000",
        "00001000",
        "00010000",
        "00010000",
        "00011000",
        "00000000",
        "10101010",
        "01010101",
        "10101010",
        "01010101",
        "10101010",
        "01010101",
        "10101010",
        "01010101"
    );
begin

    fetch_line_process: process (clk) begin
		if rising_edge(clk) then
			-- Read from Rom
			douta <= rom(to_integer(unsigned(addra)));
		end if;
	end process;

end architecture;